//
// (c) Meta Platforms, Inc. and affiliates. Confidential and proprietary.
// NOTICE OF CONFIDENTIAL AND PROPRIETARY INFORMATION & TECHNOLOGY:
// The information and technology contained herein (including the accompanying
// binary code) is the confidential information of Meta Platforms, Inc. and its
// affiliates (collectively, "Meta"). It is protected by applicable copyright
// and trade secret law, and may be claimed in one or more U.S. or foreign
// patents or pending patent applications. Meta retains all right, title and
// interest (including all intellectual property rights) in such information 
// and technology, and no licenses are hereby granted by Meta. Unauthorized
// use, reproduction, or dissemination is a violation of Meta's rights and
// is strictly prohibited.
//
// @generated
//
//------------------------------------------------------------------------------
// PACKAGE: xrbase_alfred_reg_pkg
//------------------------------------------------------------------------------
`include "uvm_macros.svh"
package xrbase_alfred_reg_pkg;
    import uvm_pkg::*;
    import fast_uvm_reg_pkg::*;
    
    `include "xrbase_alfred_reg.sv"
endpackage : xrbase_alfred_reg_pkg
