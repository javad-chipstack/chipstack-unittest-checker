//
// (c) Meta Platforms, Inc. and affiliates. Confidential and proprietary.
// NOTICE OF CONFIDENTIAL AND PROPRIETARY INFORMATION & TECHNOLOGY:
// The information and technology contained herein (including the accompanying
// binary code) is the confidential information of Meta Platforms, Inc. and its
// affiliates (collectively, "Meta"). It is protected by applicable copyright
// and trade secret law, and may be claimed in one or more U.S. or foreign
// patents or pending patent applications. Meta retains all right, title and
// interest (including all intellectual property rights) in such information 
// and technology, and no licenses are hereby granted by Meta. Unauthorized
// use, reproduction, or dissemination is a violation of Meta's rights and
// is strictly prohibited.
//
// @generated
//
// soccomp Version 10.3.0 (2ed27f84a)
// (c) Meta Platforms, Inc. and affiliates. Confidential and proprietary.
// Started soccomp on: Tue Dec 13 16:10:20 2022
// SONICS_PATH = :/nfs/project/ipgen/src/valerioc/fbrepo/common/build_root/install/studio/../extensions/include
// PYTHONPATH = PythonPathUnset
// /nfs/regress_03_ash/sonics/nightly/sonics-no-sysc-py3-daily-20221213_140241/install/studio-10.3/sonics_code/soccomp.py --relative --uvm_test --designdir ./smp --instance xrbase --post_process /nfs/project/ipgen/src/valerioc/fbrepo/common/src/neev/ipBuilder/neev/ipBuilder/GenerateIPDefs.py{"levels":"1|tile"} xrbase_alfred_smp.conf
// @generated

////////////////////////////////////////////////////////////////////////////////
// regmodel0_regmodel - Register Module Interface Definitions

interface regmodel0_regmodel_interface (
        // Interface Ports
        input                                               clk_i,
                input                                               sys_reset_ni,
                input                                               sys_test_mode_cgm_i,
                input                                               sys_test_mode_async_i,
                regmodel0_regmodel_ocp2_interface                   regmodel0_regmodel_ocp2_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src0_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src1_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src2_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src3_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src4_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src5_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src6_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src7_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src8_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src9_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src10_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src11_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src12_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src13_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src14_if,
                regmodel0_regmodel_sfdbs0_sfdb0_src_interface       regmodel0_regmodel_sfdbs0_sfdb0_src15_if,
                regmodel0_regmodel_sfdbs0_sfdb0_tgt_interface       regmodel0_regmodel_sfdbs0_sfdb0_tgt_if,
                regmodel0_regmodel_sfdbs0_ipc_sc_interface          regmodel0_regmodel_sfdbs0_ipc_sc_if,
                regmodel0_regmodel_sfdbs0_error_err_log_interface   regmodel0_regmodel_sfdbs0_error_err_log_if,
                regmodel0_regmodel_sfdbs0_error_err_data_interface  regmodel0_regmodel_sfdbs0_error_err_data_if,
                regmodel0_regmodel_sfdbs0_error_err_idx_interface   regmodel0_regmodel_sfdbs0_error_err_idx_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src0_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src1_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src2_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src3_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src4_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src5_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src6_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src7_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src8_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src9_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src10_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src11_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src12_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src13_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src14_if,
                regmodel0_regmodel_sfdbs0_sfdb1_src_interface       regmodel0_regmodel_sfdbs0_sfdb1_src15_if,
                regmodel0_regmodel_sfdbs0_sfdb1_tgt_interface       regmodel0_regmodel_sfdbs0_sfdb1_tgt_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell0_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell1_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell2_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell3_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell4_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell5_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell6_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell7_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell8_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell9_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell10_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell11_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell12_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell13_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell14_if,
                regmodel0_regmodel_fdbs0_fdb0_bell_interface        regmodel0_regmodel_fdbs0_fdb0_bell15_if,
                regmodel0_regmodel_fdbs0_fdb0_control_interface     regmodel0_regmodel_fdbs0_fdb0_control_if,
                regmodel0_regmodel_fdbs0_fdb0_enable_interface      regmodel0_regmodel_fdbs0_fdb0_enable_if,
                regmodel0_regmodel_fdbs0_fdb0_status_interface      regmodel0_regmodel_fdbs0_fdb0_status_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data0_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data1_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data2_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data3_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data4_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data5_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data6_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data7_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data8_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data9_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data10_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data11_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data12_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data13_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data14_fifo_if,
                regmodel0_regmodel_fdbs0_fdb0_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb0_data15_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell0_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell1_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell2_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell3_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell4_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell5_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell6_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell7_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell8_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell9_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell10_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell11_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell12_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell13_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell14_if,
                regmodel0_regmodel_fdbs0_fdb1_bell_interface        regmodel0_regmodel_fdbs0_fdb1_bell15_if,
                regmodel0_regmodel_fdbs0_fdb1_control_interface     regmodel0_regmodel_fdbs0_fdb1_control_if,
                regmodel0_regmodel_fdbs0_fdb1_enable_interface      regmodel0_regmodel_fdbs0_fdb1_enable_if,
                regmodel0_regmodel_fdbs0_fdb1_status_interface      regmodel0_regmodel_fdbs0_fdb1_status_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data0_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data1_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data2_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data3_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data4_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data5_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data6_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data7_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data8_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data9_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data10_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data11_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data12_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data13_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data14_fifo_if,
                regmodel0_regmodel_fdbs0_fdb1_data_fifo_interface   regmodel0_regmodel_fdbs0_fdb1_data15_fifo_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner0_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner1_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner2_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner3_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner4_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner5_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner6_if,
                regmodel0_regmodel_smutex0_owner_interface          regmodel0_regmodel_smutex0_owner7_if,
                regmodel0_regmodel_smutex0_ipc_sc_interface         regmodel0_regmodel_smutex0_ipc_sc_if,
                regmodel0_regmodel_smutex0_timeout_interface        regmodel0_regmodel_smutex0_timeout_if,
                regmodel0_regmodel_smutex0_error_err_log_interface  regmodel0_regmodel_smutex0_error_err_log_if,
                regmodel0_regmodel_smutex0_error_err_data_interface regmodel0_regmodel_smutex0_error_err_data_if,
                regmodel0_regmodel_smutex0_error_err_idx_interface  regmodel0_regmodel_smutex0_error_err_idx_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex0_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex1_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex2_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex3_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex4_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex5_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex6_if,
                regmodel0_regmodel_mutex0_mutex_interface           regmodel0_regmodel_mutex0_mutex7_if,
                regmodel0_regmodel_web0_control_interface           regmodel0_regmodel_web0_control_if,
                regmodel0_regmodel_web0_event_interface             regmodel0_regmodel_web0_event_if,
                regmodel0_regmodel_web0_wake_enable0_interface      regmodel0_regmodel_web0_wake_enable0_if,
                regmodel0_regmodel_web0_wake_enable1_interface      regmodel0_regmodel_web0_wake_enable1_if,
                regmodel0_regmodel_web0_input_invert0_interface     regmodel0_regmodel_web0_input_invert0_if,
                regmodel0_regmodel_web0_input_invert1_interface     regmodel0_regmodel_web0_input_invert1_if,
                regmodel0_regmodel_web1_control_interface           regmodel0_regmodel_web1_control_if,
                regmodel0_regmodel_web1_event_interface             regmodel0_regmodel_web1_event_if,
                regmodel0_regmodel_web1_wake_enable0_interface      regmodel0_regmodel_web1_wake_enable0_if,
                regmodel0_regmodel_web1_wake_enable1_interface      regmodel0_regmodel_web1_wake_enable1_if,
                regmodel0_regmodel_web1_input_invert0_interface     regmodel0_regmodel_web1_input_invert0_if,
                regmodel0_regmodel_web1_input_invert1_interface     regmodel0_regmodel_web1_input_invert1_if    
    );
endinterface

